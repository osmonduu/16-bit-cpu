`define READ 0
`define WRITE 1
`define PCR 16 // program counter index
`define tick #1clock=1;#1clock=0
`define dbg